library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

ENTITY FRAME_BUFFER IS
	PORT(
		-- IN SIGNALS
		RD_VALID: IN STD_LOGIC;
		RD_DATA: IN STD_LOGIC_VECTOR(7 downto 0);
		
		--SRAM
		SRAM_CE_N, SRAM_OE_N, SRAM_WE_N, SRAM_UB_N, SRAM_LB_N: OUT STD_LOGIC;
		SRAM_ADDR: OUT STD_LOGIC_VECTOR(17 downto 0);
		SRAM_DQ: INOUT STD_LOGIC_VECTOR(15 downto 0);
		
		-- OUT SIGNALS
		WR_FULL: IN STD_LOGIC;
		WR_REQ: OUT STD_LOGIC;
		WR_DATA: OUT STD_LOGIC_VECTOR(7 downto 0);
		
		--CLOCK AND RESET
		CLK, RESET: IN STD_LOGIC
	);
END FRAME_BUFFER;

ARCHITECTURE FRAME_BUFFER_ARCH OF FRAME_BUFFER IS
	--BETWEEN WRITER AND CONTROLLER
	SIGNAL WR_ACK_REG, WR_REQ_REG: STD_LOGIC;
	SIGNAL WR_DATA_REG: STD_LOGIC_VECTOR(15 DOWNTO 0);
	SIGNAL WR_ADDR_REG: STD_LOGIC_VECTOR(17 DOWNTO 0);
	
	--BETWEEN READER AND CONTROLLER
	SIGNAL RD_REQ_REG: STD_LOGIC;
	SIGNAL RD_ACK_REG: STD_LOGIC;
	SIGNAL RD_ADDR_REG: STD_LOGIC_VECTOR(17 downto 0);
	SIGNAL RD_DATA_REG: STD_LOGIC_VECTOR(15 downto 0);
	
	COMPONENT SRAM_WRITER IS
		PORT(
			-- FIFO CHANNEL --
			RD_VALID: IN STD_LOGIC;
			RD_DATA: IN STD_LOGIC_VECTOR(7 downto 0);
			
			-- SRAM CONTROLLER CHANNEL --
			WR_ACK : IN STD_LOGIC;
			DATA_OUT: OUT STD_LOGIC_VECTOR(15 downto 0);
			WR_ADDR : OUT STD_LOGIC_VECTOR(17 downto 0);
			WR      : OUT STD_LOGIC;
			
			-- CLK and RESET --
			CLK, RESET: IN STD_LOGIC			
		);
	END COMPONENT SRAM_WRITER;
	
	COMPONENT SRAM_CONTROLLER IS
	PORT(
		-- READ CHANNEL --
		RD_REQ: IN STD_LOGIC;
		RD_ACK: OUT STD_LOGIC;
		RD_ADDR: IN STD_LOGIC_VECTOR(17 downto 0);
		RD_DATA: OUT STD_LOGIC_VECTOR(15 downto 0);
		
		-- WRITE CHANNEL --
		WR_REQ: IN STD_LOGIC;
		WR_ACK: OUT STD_LOGIC;
		WR_ADDR: IN STD_LOGIC_VECTOR(17 downto 0);
		WR_DATA: IN STD_LOGIC_VECTOR(15 downto 0);
		
		-- SRAM BUS SIGNALS --
		SRAM_CE_N, SRAM_OE_N, SRAM_WE_N, SRAM_UB_N, SRAM_LB_N: OUT STD_LOGIC;
		SRAM_ADDR: OUT STD_LOGIC_VECTOR(17 downto 0);
		SRAM_DQ: INOUT STD_LOGIC_VECTOR(15 downto 0);
		
		-- CLK and RESET --
		CLK, RESET: IN STD_LOGIC	
	);
	END COMPONENT SRAM_CONTROLLER;
	
	COMPONENT SRAM_READER IS
	PORT(
		-- FIFO CHANNEL --
		WR_FULL: IN STD_LOGIC;
		WR_REQ: OUT STD_LOGIC;
		WR_DATA: OUT STD_LOGIC_VECTOR(7 downto 0);
		
		-- SRAM CONTROLLER CHANNEL --
		RD_ACK: IN STD_LOGIC;
		DATA_IN: IN STD_LOGIC_VECTOR(15 downto 0);
		RD_ADDR: OUT STD_LOGIC_VECTOR(17 downto 0);
		RD: OUT STD_LOGIC;
		
		-- CLK and RESET --
		CLK, RESET: IN STD_LOGIC
	);
	END COMPONENT SRAM_READER;
	
 BEGIN
	WRITER: SRAM_WRITER PORT MAP(RD_VALID, RD_DATA, WR_ACK_REG, WR_DATA_REG, WR_ADDR_REG, WR_REQ_REG, CLK, RESET);
	CONTROLLER: SRAM_CONTROLLER PORT MAP(
		RD_REQ_REG, RD_ACK_REG, RD_ADDR_REG, RD_DATA_REG,
		WR_REQ_REG, WR_ACK_REG, WR_ADDR_REG,WR_DATA_REG,
		SRAM_CE_N, SRAM_OE_N, SRAM_WE_N, SRAM_UB_N, SRAM_LB_N, SRAM_ADDR,SRAM_DQ,
		CLK, RESET
	);
	READER: SRAM_READER PORT MAP(WR_FULL, WR_REQ, WR_DATA, RD_ACK_REG, RD_DATA_REG, RD_ADDR_REG, RD_REQ_REG, CLK, RESET);
 END FRAME_BUFFER_ARCH;
