library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

ENTITY VGA_CONTROLLER IS
PORT(

	HSYNC: OUT STD_LOGIC;
	VSYNC: OUT STD_LOGIC;
	R: OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
	G: OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
	B: OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
	R_IN: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
	G_IN: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
	B_IN: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
	DATA_ACK: OUT STD_LOGIC;
	
	CLK: IN STD_LOGIC;
	RST: IN STD_LOGIC
);
END VGA_CONTROLLER;


ARCHITECTURE VGA_CONTROLLER_ARCH OF VGA_CONTROLLER IS
	--640x480 @ 60 Hz pixel clock 25.175MHz
	
	CONSTANT HOR: INTEGER := 640;
	CONSTANT HORIZONTAL_FP: INTEGER := 16;
	CONSTANT HORIZONTAL_BP: INTEGER := 48;
	CONSTANT HORIZONTAL_SYNC_PULSE: INTEGER := 96;
	
	CONSTANT H_STARTSYNC: INTEGER := HOR + HORIZONTAL_FP;
	CONSTANT H_ENDSYNC: INTEGER := H_STARTSYNC + HORIZONTAL_SYNC_PULSE;
	CONSTANT HOR_TOT: INTEGER := HOR + HORIZONTAL_BP + HORIZONTAL_FP + HORIZONTAL_SYNC_PULSE;
	
	CONSTANT VER: INTEGER := 480;
	CONSTANT VERTICAL_FP: INTEGER := 10;
	CONSTANT VERTICAL_BP: INTEGER := 33;
	CONSTANT VERTICAL_SYNC_PULSE: INTEGER := 2;
	
	CONSTANT V_STARTSYNC: INTEGER := VER + VERTICAL_FP;
	CONSTANT V_ENDSYNC: INTEGER := V_STARTSYNC + VERTICAL_SYNC_PULSE;
	CONSTANT VER_TOT: INTEGER := VER + VERTICAL_BP + VERTICAL_FP + VERTICAL_SYNC_PULSE;
	
	SIGNAL BLANK: STD_LOGIC := '1';
	BEGIN

	PROCESS(CLK, RST)
	VARIABLE HPOS: INTEGER RANGE 0 TO HOR_TOT-1:=0;
	VARIABLE VPOS: INTEGER RANGE 0 TO VER_TOT-1:=0;
		BEGIN
			IF(RST = '1')
			THEN
				HPOS := 0;
				VPOS := 0;
				BLANK <= '1';
				R<=(others=>'0');
				G<=(others=>'0');
				B<=(others=>'0');
				
			ELSIF(RISING_EDGE(CLK))
			THEN
				--AGGIORNAMENTO POSIZIONE
				IF(HPOS = HOR_TOT-1)
				THEN
					HPOS := 0;
					VPOS := (VPOS + 1) MOD VER_TOT;
				ELSE
					HPOS := HPOS+1;
				END IF;
				--FINE AGGIORNAMENTO
				
				--GESTIONE FLUSSO OUTPUT
				IF(BLANK = '1')
				THEN
					R<=(others=>'0');
					G<=(others=>'0');
					B<=(others=>'0');
				ELSE
					R <= R_IN;
					G <= G_IN;
					B <= B_IN;
				END IF;
				--FINE GESTIONE FLUSSO OUTPUT
				
				--BLANK TIMING
				IF(VPOS >=  VER)
				THEN
					BLANK <= '1';
					ELSE
					IF(HPOS < HOR)
					THEN
						BLANK <='0';
					ELSE
						BLANK <='1';
					END IF;					
				END IF;
				--FINE BLANK TIMING
				
				-- SYNC TIMING
				IF(HPOS > H_STARTSYNC AND HPOS <= H_ENDSYNC)
				THEN
					HSYNC <= '0';
				ELSE
					HSYNC <= '1';
				END IF;
				
				IF(VPOS >= V_STARTSYNC AND VPOS < V_ENDSYNC)
				THEN
					VSYNC <= '0';
				ELSE
					VSYNC <= '1';
				END IF;
				-- FINE SYNC TIMING
			END IF;
		END PROCESS;
		
		--LOGICA NEGATA
		DATA_ACK <= NOT BLANK;
	 
 END VGA_CONTROLLER_ARCH;